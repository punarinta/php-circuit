V1 0 UCC DC 1
R1 UCC A 5
C1 A 0 100n

.TRAN 50n 500n
.PLOT TRAN V(A)
